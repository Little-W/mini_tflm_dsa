`timescale 1ns / 1ps

module tb_compute_core;
    localparam int unsigned SIZE = 4;
    localparam int unsigned DATA_WIDTH = 16;

    // 添加 ANSI 颜色常量
    localparam string C_GREEN = "\033[0;32m";
    localparam string C_RED   = "\033[0;31m";
    localparam string C_RESET = "\033[0m";

    // clock
    logic clk;
    initial clk = 0;
    always #5 clk <= ~clk;  // 100MHz

    // Instantiate interface
    tb_compute_core_if tb_if(clk);

    // memories for stimuli and expected
    // 先用原始位宽的临时数组读文件，再打包到32位数组
    logic signed [           7:0] weight_mem_raw        [  SIZE*16];  // 64B
    logic signed [DATA_WIDTH-1:0] ia_mem_raw            [  SIZE*16];  // 64 halfwords
    localparam int WeightWords = (SIZE*16)/4;  // 64B / 4 = 16
    localparam int IaWords     = (SIZE*16)/2;  // 64H / 2 = 32
    logic        [          31:0] weight_mem            [WeightWords];
    logic        [          31:0] ia_mem                [  IaWords];
    logic signed [          31:0] exp_mem               [SIZE*SIZE];  // SIZE x SIZE
    // 新增：每个输出通道的32位偏置
    logic signed [          31:0] bias_mem              [     SIZE];

    // capture buffer
    logic signed [          31:0] out_buf               [SIZE*SIZE];
    integer                       out_rows;

    // helpers
    integer                       errors;
    integer                       idx;
    integer                       NUM_K;
    integer                       NUM_SEG;

    // tile_buf声明移到模块顶部
    logic signed [7:0] tile_buf [SIZE][SIZE];

    // init defaults
    initial begin
        out_rows             = 0;
        errors               = 0;
        NUM_K                = 16;
        NUM_SEG              = NUM_K / SIZE;
    end

    // DUT
    compute_core #(
        .SIZE      (SIZE),
        .DATA_WIDTH(DATA_WIDTH)
    ) u_dut (
        .clk                  (clk),
        .store_weight_req     (tb_if.store_weight_req),
        .weight_in            (tb_if.weight_in),
        .ia_vec_in            (tb_if.ia_vec_in),
        .ia_row_valid         (tb_if.ia_row_valid),
        .ia_calc_done         (tb_if.ia_calc_done),
        .ia_is_init_data      (tb_if.ia_is_init_data),
        .bias_in              (tb_if.bias_in),
        .acc_data_out         (tb_if.acc_data_out),
        .acc_data_valid       (tb_if.acc_data_valid),
        .tile_calc_over       (tb_if.tile_calc_over),
        .partial_sum_calc_over(tb_if.partial_sum_calc_over)
    );

    // waveform dump
    initial begin
        $dumpfile("wave.vcd");
        $dumpvars(0, tb_compute_core);
    end

    // capture outputs when valid: each cycle a row of SIZE outputs
    always @(posedge clk) begin
        if (tb_if.acc_data_valid) begin
            for (int c = 0; c < SIZE; c++) begin
                out_buf[out_rows*SIZE+c] <= tb_if.acc_data_out[c];
            end
            out_rows <= out_rows + 1;
        end
    end

    // main stimulus
    initial begin
        // load data from files generated by Python（先读原始位宽临时数组）
        $readmemh("/home/etc/FPGA/tflm_ai_dsa/test/compute_core/weight_mem.hex", weight_mem_raw);
        $readmemh("/home/etc/FPGA/tflm_ai_dsa/test/compute_core/ia_mem.hex", ia_mem_raw);
        $readmemh("/home/etc/FPGA/tflm_ai_dsa/test/compute_core/expected_out.hex", exp_mem);
        // 读取偏置
        $readmemh("/home/etc/FPGA/tflm_ai_dsa/test/compute_core/bias_mem.hex", bias_mem);

        // 将临时数组打包到32位数组：权重4x8bit/word，IA 2x16bit/word
        for (int i = 0; i < WeightWords; i++) begin
            weight_mem[i][7:0]    = weight_mem_raw[i*4+0];
            weight_mem[i][15:8]   = weight_mem_raw[i*4+1];
            weight_mem[i][23:16]  = weight_mem_raw[i*4+2];
            weight_mem[i][31:24]  = weight_mem_raw[i*4+3];
        end
        for (int i = 0; i < IaWords; i++) begin
            ia_mem[i][15:0]  = ia_mem_raw[i*2+0];
            ia_mem[i][31:16] = ia_mem_raw[i*2+1];
        end

        // small delay for stability
        repeat (5) @(tb_if.cb);

        // 分段（K方向按SIZE=4切分）：每段先加载4行权重，再输入4拍IA
        for (int seg = 0; seg < NUM_SEG; seg++) begin
            // 在加载下一段权重前，必须等待上一段部分和完成
            if (seg != 0) begin
                $display("[TB] Wait partial_sum_calc_over before next weight seg=%0d", seg);
                wait (tb_if.partial_sum_calc_over == 1'b1);
                @(tb_if.cb);
            end

            // 1) 加载本段权重：store_weight_req=1，每拍一行（共SIZE行）
            $display("[TB] Loading weight tile seg=%0d", seg);
            load_weight_tile(seg);

            // 加载对应通道偏置（仅首段加载，否则清零）
            load_bias(seg);

            // 空转一拍，便于DUT内部状态稳定
            @(tb_if.cb);

            // 2) 输入本段IA向量：ia_row_valid=1，连续SIZE拍
            $display("[TB] Streaming IA tile seg=%0d", seg);
            stream_ia_tile(seg);
        end

        // 3) 等待整个tile完成，再进行结果对比
        $display("[TB] Waiting for tile_calc_over...");
        wait (tb_if.tile_calc_over == 1'b1);
        $display("[TB] tile_calc_over detected");
        repeat (2) @(tb_if.cb);

        if (out_rows < SIZE) begin
            $display("ERROR: output rows=%0d < expected=%0d", out_rows, SIZE);
            errors = errors + 1;
        end
        for (int r = 0; r < SIZE; r++) begin
            for (int c = 0; c < SIZE; c++) begin
                idx = r * SIZE + c;
                if (out_buf[idx] !== exp_mem[idx]) begin
                    $display("MISMATCH r=%0d c=%0d", r, c);
                    $display("  got=%0d (0x%08h)", out_buf[idx], out_buf[idx]);
                    $display("  exp=%0d (0x%08h)", exp_mem[idx], exp_mem[idx]);
                    errors = errors + 1;
                end
            end
        end

        if (errors == 0) $display("%sPASS: compute_core 4x16 * 16x4 matched expected%s", C_GREEN, C_RESET);
        else               $display("%sFAIL: %0d mismatches%s", C_RED, errors, C_RESET);

        #20;
        $finish;
    end

    // 偏置加载任务。仅在首个seg加载偏置，其余seg清零。
    task automatic load_bias(input int seg);
        begin
            if (seg == 0) begin
                for (int c = 0; c < SIZE; c++) begin
                    tb_if.cb.bias_in[c] <= bias_mem[c];
                end
            end else begin
                for (int c = 0; c < SIZE; c++) begin
                    tb_if.cb.bias_in[c] <= 32'sd0;
                end
            end
        end
    endtask

    task automatic load_weight_tile(input int seg);
        begin
            tb_if.cb.store_weight_req <= 1'b1;
            // 每列一次性读取4个8bit权重（一个32bit）
            for (int c = 0; c < SIZE; c++) begin
                int base_idx8;
                logic [31:0] w32;
                base_idx8 = (seg * SIZE) + c * NUM_K; // 对齐到4字节
                w32       = weight_mem[base_idx8 >> 2];
                // 展开为4个字节，避免动态部分选择
                tile_buf[0][c] = $signed(w32[7:0]);
                tile_buf[1][c] = $signed(w32[15:8]);
                tile_buf[2][c] = $signed(w32[23:16]);
                tile_buf[3][c] = $signed(w32[31:24]);
            end
            // 按行输出
            for (int k = SIZE - 1; k >= 0; k--) begin
                for (int j = 0; j < SIZE; j++) begin
                    tb_if.cb.weight_in[j] <= tile_buf[k][j];
                end
                @(tb_if.cb);
            end
            tb_if.cb.store_weight_req <= 1'b0;
        end
    endtask

    task automatic stream_ia_tile(input int seg);
        begin
            tb_if.cb.ia_row_valid <= 1'b1;
            tb_if.cb.ia_is_init_data <= (seg == 0);
            tb_if.cb.ia_calc_done <= (seg == (NUM_SEG - 1));
            for (int k = 0; k < SIZE; k++) begin
                int base16;
                logic [31:0] p0, p1;
                base16 = seg * SIZE + k * NUM_K; // 对齐到2个16bit
                p0 = ia_mem[ base16       >> 1]; // 包含base16, base16+1
                p1 = ia_mem[(base16 + 2) >> 1]; // 包含base16+2, base16+3
                tb_if.cb.ia_vec_in[0] <= p0[15:0];
                tb_if.cb.ia_vec_in[1] <= p0[31:16];
                tb_if.cb.ia_vec_in[2] <= p1[15:0];
                tb_if.cb.ia_vec_in[3] <= p1[31:16];
                @(tb_if.cb);
            end
            tb_if.cb.ia_row_valid <= 1'b0;
            tb_if.cb.ia_is_init_data <= 1'b0;
            tb_if.cb.ia_calc_done <= 1'b0;
            for (int r = 0; r < SIZE; r++) tb_if.cb.ia_vec_in[r] <= 0;
        end
    endtask

endmodule
