`include "define.svh"
module global_controller #(
) (
);

endmodule